module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 ;
  output y0 ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n8 = x1 | x2 ;
  assign n9 = x1 & x2 ;
  assign n10 = x0 | n9 ;
  assign n11 = n8 | n10 ;
  assign n12 = x3 | x4 ;
  assign n13 = x5 & x6 ;
  assign n14 = n12 & n13 ;
  assign n15 = x3 & x4 ;
  assign n16 = x5 | x6 ;
  assign n17 = n15 & n16 ;
  assign n18 = n14 | n17 ;
  assign n19 = n11 & n18 ;
  assign n20 = x0 & n9 ;
  assign n21 = n12 | n13 ;
  assign n22 = n15 | n16 ;
  assign n23 = n21 | n22 ;
  assign n24 = n20 & n23 ;
  assign n25 = n19 | n24 ;
  assign n26 = n14 & n17 ;
  assign n27 = n8 & n10 ;
  assign n28 = n21 & n22 ;
  assign n29 = n27 & n28 ;
  assign n30 = n26 | n29 ;
  assign n31 = n25 | n30 ;
  assign y0 = n31 ;
endmodule
